`include "TIME_SCALE.svh"
`include "SAL_DDR_PARAMS.svh"

module SAL_DDR_CTRL
(
    // clock & reset
    input                       clk,
    input                       rst_n,

    // APB interface
    APB_IF.SLV                  apb_if,

    // AXI interface
    AXI_IF.SLV                  axi_if,

    // DFI interface
    DFI_CTRL_IF.SRC             dfi_ctrl_if,
    DFI_WR_IF.SRC               dfi_wr_if,
    DFI_RD_IF.DST               dfi_rd_if
);

    // timing parameters
    TIMING_IF                   timing_if();

    // requests to a bank
    REQ_IF                      bk_req_if_arr[`DRAM_BK_CNT](.clk(clk), .rst_n(rst_n));
    // requests to the scheduler
    SCHED_IF                    bk_sched_if_arr[`DRAM_BK_CNT] ();
    // scheduling output
    SCHED_IF                    sched_if();

    AXI_IF                      axi_internal_if     (.clk(clk), .rst_n(rst_n));

    // Configurations
    SAL_CFG                         u_cfg
    (
        .clk                        (clk),
        .rst_n                      (rst_n),

        .apb_if                     (apb_if),

        .timing_if                  (timing_if)
    );

    SAL_WR_CTRL                     u_wr_ctrl
    (
        .clk                        (clk),
        .rst_n                      (rst_n),

        .timing_if                  (timing_if),
        .sched_if                   (sched_if),

        .axi_aw_if                  (axi_if),
        .axi_w_if                   (axi_if),
        .axi_b_if                   (axi_if),

        .axi_aw2_if                 (axi_internal_if),
        .dfi_wr_if                  (dfi_wr_if)
    );

    SAL_ADDR_DECODER                u_decoder
    (
        .clk                        (clk),
        .rst_n                      (rst_n),

        .axi_ar_if                  (axi_if.SLV_AR),
        .axi_aw_if                  (axi_internal_if),

        .req_if_arr                 (bk_req_if_arr)
    );

    genvar geni;

    generate
        for (geni=0; geni<`DRAM_BK_CNT; geni=geni+1) begin  : BK
            SAL_BK_CTRL                     u_bank_ctrl
            (
                .clk                        (clk),
                .rst_n                      (rst_n),
        
                .timing_if                  (timing_if),
        
                .req_if                     (bk_req_if_arr[geni]),
                .sched_if                   (bk_sched_if_arr[geni]),
        
                .ref_req_i                  (1'b0),
                .ref_gnt_o                  ()
            );
        end
    endgenerate

    SAL_SCHED                       u_sched
    (
        .clk                        (clk),
        .rst_n                      (rst_n),

        .bk_sched_if_arr            (bk_sched_if_arr),
        .sched_if                   (sched_if)
    );

    SAL_CTRL_ENCODER                u_encoder
    (
        .clk                        (clk),
        .rst_n                      (rst_n),

        .sched_if                   (sched_if),
        .dfi_ctrl_if                (dfi_ctrl_if)
    );

    SAL_RD_CTRL                     u_rd_ctrl
    (
        .clk                        (clk),
        .rst_n                      (rst_n),

        .timing_if                  (timing_if),
        .sched_if                   (sched_if),
        .dfi_rd_if                  (dfi_rd_if),
        .axi_r_if                   (axi_if)
    );

endmodule // SAL_DDR_CTRL
